//=================================================================
// Class Description: Data items for APB UVC
// Project Name:	    renas mcu
// Ho Chi Minh University of Technology
// Email: 			quanghungbk1999@gmail.com  
// Version  Date        Author    Description
// v0.0     18.03.2021  hungbk99  First Creation  
//=================================================================

typedef enum bit {APB_READ, APB_WRITE} apb_direction_enum;
